module alu8bit(opcode,in1,in2,result,flagc,flagz);
input [7:0]in1,in2;
input [2:0]opcode;
output reg [15:0] result = 16'b0;
output reg flagz=1'b0;
output reg flagc=1'b0;
parameter [2:0] ADD =3'b000,
SUB=3'b001,MUL=3'b010,AND=3'b011,
OR=3'b100,NAND=3'b101,NOR=3'b110,
XOR=3'b111;
always@(opcode,in1,in2)
begin
case(opcode)
ADD: begin 
result =in1+in2;
flagc=result[8];
flagz=(result==16'b0);
end

SUB: begin
result=in1-in2;
flagc=result[8];
flagz=(result==16'b0);
end

MUL: begin
result=in1*in2;
flagz=(result==16'b0);
end

AND: begin
result=in1&in2;
flagz=(result==16'b0);
end


OR: begin
result=in1|in2;
flagz=(result==16'b0);
end


NAND: begin
result=~(in1&in2);
flagz=(result==16'b0);
end


NOR: begin
result=~(in1|in2);
flagz=(result==16'b0);
end

XOR: begin
result=(in1^in2);
flagz=(result==16'b0);
end
endcase
end
endmodule
